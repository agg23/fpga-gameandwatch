// Build ID Verilog Module
`define BUILD_DATE "20230622"
`define BUILD_HASH "afc5696b"
