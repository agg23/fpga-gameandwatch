// Build ID Verilog Module
`define BUILD_DATE "20230624"
`define BUILD_HASH "39c3a75e"
