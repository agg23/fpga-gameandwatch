// Build ID Verilog Module
`define BUILD_DATE "20230626"
`define BUILD_HASH "3d8d9c4a"
