//------------------------------------------------------------------------------
// SPDX-License-Identifier: MIT
// SPDX-FileType: SOURCE
// SPDX-FileCopyrightText: (c) 2023, agg23
//------------------------------------------------------------------------------

`default_nettype none

module gameandwatch ();

endmodule
