// Build ID Verilog Module
`define BUILD_DATE "20230623"
`define BUILD_HASH "02d09629"
